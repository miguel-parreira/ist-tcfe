.OP
R1 v1 v2 1.02815650737k
R2 v3 v2 2.07414279923k
R3 v2 v5 3.06367122238k
R4 v5 GND 4.06922855851k
R5 v5 v6 3.03804085665k
R6 GND v7 2.05484565321k
R7 vaux v8 1.02936604691k
Vs v1 GND 0
vamp v7 vaux 0
hVc  v5 v8  vamp  8.1158893784k
gVc v6 v3 v2 v5 7.2545889117m
.END

